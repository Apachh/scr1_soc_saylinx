module saylinx_scr1 (

);